interface adder_if;

    logic [2:0] a;
    logic [2:0] b;
    logic cin;
    logic [3:0] dout;

endinterface